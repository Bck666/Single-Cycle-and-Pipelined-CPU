module InstructionMemory(
	input      [32 -1:0] Address, 
	output reg [32 -1:0] Instruction
);
	
	always @(*)
		case (Address[13:2])

			// -------- Paste Binary Instruction Below (Inst-q1.txt, Inst-q2.txt, Inst-q3.txt)
10'd0:  Instruction <= 32'h24080000;
            10'd1:  Instruction <= 32'h8d100000;
            10'd2:  Instruction <= 32'h00102021;
            10'd3:  Instruction <= 32'h21050004;
            10'd4:  Instruction <= 32'h0c100142;
            10'd5:  Instruction <= 32'h24080001;
            10'd6:  Instruction <= 32'h24091068;
            10'd7:  Instruction <= 32'h240b0000;
            10'd8:  Instruction <= 32'h21290004;
            10'd9:  Instruction <= 32'h8d240000;
            10'd10:  Instruction <= 32'h01645820;
            10'd11:  Instruction <= 32'h21080001;
            10'd12:  Instruction <= 32'h0110082a;
            10'd13:  Instruction <= 32'h1420fffa;
            10'd14:  Instruction <= 32'h0010c880;
            10'd15:  Instruction <= 32'h232a1068;
            10'd16:  Instruction <= 32'had4b0000;
            10'd17:  Instruction <= 32'h3c014000;
            10'd18:  Instruction <= 32'h34340010;
            10'd19:  Instruction <= 32'hae800000;
            10'd20:  Instruction <= 32'h8d480000;
            10'd21:  Instruction <= 32'h00082700;
            10'd22:  Instruction <= 32'h00042702;
            10'd23:  Instruction <= 32'h24090000;
            10'd24:  Instruction <= 32'h1089001e;
            10'd25:  Instruction <= 32'h24090001;
            10'd26:  Instruction <= 32'h1089001e;
            10'd27:  Instruction <= 32'h24090002;
            10'd28:  Instruction <= 32'h1089001e;
            10'd29:  Instruction <= 32'h24090003;
            10'd30:  Instruction <= 32'h1089001e;
            10'd31:  Instruction <= 32'h24090004;
            10'd32:  Instruction <= 32'h1089001e;
            10'd33:  Instruction <= 32'h24090005;
            10'd34:  Instruction <= 32'h1089001e;
            10'd35:  Instruction <= 32'h24090006;
            10'd36:  Instruction <= 32'h1089001e;
            10'd37:  Instruction <= 32'h24090007;
            10'd38:  Instruction <= 32'h1089001e;
            10'd39:  Instruction <= 32'h24090008;
            10'd40:  Instruction <= 32'h1089001e;
            10'd41:  Instruction <= 32'h24090009;
            10'd42:  Instruction <= 32'h1089001e;
            10'd43:  Instruction <= 32'h2409000a;
            10'd44:  Instruction <= 32'h1089001e;
            10'd45:  Instruction <= 32'h2409000b;
            10'd46:  Instruction <= 32'h1089001e;
            10'd47:  Instruction <= 32'h2409000c;
            10'd48:  Instruction <= 32'h1089001e;
            10'd49:  Instruction <= 32'h2409000d;
            10'd50:  Instruction <= 32'h1089001e;
            10'd51:  Instruction <= 32'h2409000e;
            10'd52:  Instruction <= 32'h1089001e;
            10'd53:  Instruction <= 32'h2409000f;
            10'd54:  Instruction <= 32'h1089001e;
            10'd55:  Instruction <= 32'h24040040;
            10'd56:  Instruction <= 32'h08100057;
            10'd57:  Instruction <= 32'h24040079;
            10'd58:  Instruction <= 32'h08100057;
            10'd59:  Instruction <= 32'h24040024;
            10'd60:  Instruction <= 32'h08100057;
            10'd61:  Instruction <= 32'h24040030;
            10'd62:  Instruction <= 32'h08100057;
            10'd63:  Instruction <= 32'h24040019;
            10'd64:  Instruction <= 32'h08100057;
            10'd65:  Instruction <= 32'h24040012;
            10'd66:  Instruction <= 32'h08100057;
            10'd67:  Instruction <= 32'h24040002;
            10'd68:  Instruction <= 32'h08100057;
            10'd69:  Instruction <= 32'h24040078;
            10'd70:  Instruction <= 32'h08100057;
            10'd71:  Instruction <= 32'h24040000;
            10'd72:  Instruction <= 32'h08100057;
            10'd73:  Instruction <= 32'h24040010;
            10'd74:  Instruction <= 32'h08100057;
            10'd75:  Instruction <= 32'h24040008;
            10'd76:  Instruction <= 32'h08100057;
            10'd77:  Instruction <= 32'h24040003;
            10'd78:  Instruction <= 32'h08100057;
            10'd79:  Instruction <= 32'h24040046;
            10'd80:  Instruction <= 32'h08100057;
            10'd81:  Instruction <= 32'h24040021;
            10'd82:  Instruction <= 32'h08100057;
            10'd83:  Instruction <= 32'h24040006;
            10'd84:  Instruction <= 32'h08100057;
            10'd85:  Instruction <= 32'h2404000e;
            10'd86:  Instruction <= 32'h08100057;
            10'd87:  Instruction <= 32'h20840e00;
            10'd88:  Instruction <= 32'h00082e00;
            10'd89:  Instruction <= 32'h00052e02;
            10'd90:  Instruction <= 32'h00052902;
            10'd91:  Instruction <= 32'h0005c021;
            10'd92:  Instruction <= 32'h24090000;
            10'd93:  Instruction <= 32'h10a9001e;
            10'd94:  Instruction <= 32'h24090001;
            10'd95:  Instruction <= 32'h10a9001e;
            10'd96:  Instruction <= 32'h24090002;
            10'd97:  Instruction <= 32'h10a9001e;
            10'd98:  Instruction <= 32'h24090003;
            10'd99:  Instruction <= 32'h10a9001e;
            10'd100:  Instruction <= 32'h24090004;
            10'd101:  Instruction <= 32'h10a9001e;
            10'd102:  Instruction <= 32'h24090005;
            10'd103:  Instruction <= 32'h10a9001e;
            10'd104:  Instruction <= 32'h24090006;
            10'd105:  Instruction <= 32'h10a9001e;
            10'd106:  Instruction <= 32'h24090007;
            10'd107:  Instruction <= 32'h10a9001e;
            10'd108:  Instruction <= 32'h24090008;
            10'd109:  Instruction <= 32'h10a9001e;
            10'd110:  Instruction <= 32'h24090009;
            10'd111:  Instruction <= 32'h10a9001e;
            10'd112:  Instruction <= 32'h2409000a;
            10'd113:  Instruction <= 32'h10a9001e;
            10'd114:  Instruction <= 32'h2409000b;
            10'd115:  Instruction <= 32'h10a9001e;
            10'd116:  Instruction <= 32'h2409000c;
            10'd117:  Instruction <= 32'h10a9001e;
            10'd118:  Instruction <= 32'h2409000d;
            10'd119:  Instruction <= 32'h10a9001e;
            10'd120:  Instruction <= 32'h2409000e;
            10'd121:  Instruction <= 32'h10a9001e;
            10'd122:  Instruction <= 32'h2409000f;
            10'd123:  Instruction <= 32'h10a9001e;
            10'd124:  Instruction <= 32'h24050040;
            10'd125:  Instruction <= 32'h0810009c;
            10'd126:  Instruction <= 32'h24050079;
            10'd127:  Instruction <= 32'h0810009c;
            10'd128:  Instruction <= 32'h24050024;
            10'd129:  Instruction <= 32'h0810009c;
            10'd130:  Instruction <= 32'h24050030;
            10'd131:  Instruction <= 32'h0810009c;
            10'd132:  Instruction <= 32'h24050019;
            10'd133:  Instruction <= 32'h0810009c;
            10'd134:  Instruction <= 32'h24050012;
            10'd135:  Instruction <= 32'h0810009c;
            10'd136:  Instruction <= 32'h24050002;
            10'd137:  Instruction <= 32'h0810009c;
            10'd138:  Instruction <= 32'h24050078;
            10'd139:  Instruction <= 32'h0810009c;
            10'd140:  Instruction <= 32'h24050000;
            10'd141:  Instruction <= 32'h0810009c;
            10'd142:  Instruction <= 32'h24050010;
            10'd143:  Instruction <= 32'h0810009c;
            10'd144:  Instruction <= 32'h24050008;
            10'd145:  Instruction <= 32'h0810009c;
            10'd146:  Instruction <= 32'h24050003;
            10'd147:  Instruction <= 32'h0810009c;
            10'd148:  Instruction <= 32'h24050046;
            10'd149:  Instruction <= 32'h0810009c;
            10'd150:  Instruction <= 32'h24050021;
            10'd151:  Instruction <= 32'h0810009c;
            10'd152:  Instruction <= 32'h24050006;
            10'd153:  Instruction <= 32'h0810009c;
            10'd154:  Instruction <= 32'h2405000e;
            10'd155:  Instruction <= 32'h0810009c;
            10'd156:  Instruction <= 32'h20a50d00;
            10'd157:  Instruction <= 32'h00083500;
            10'd158:  Instruction <= 32'h00063502;
            10'd159:  Instruction <= 32'h00063202;
            10'd160:  Instruction <= 32'h24090000;
            10'd161:  Instruction <= 32'h10c9001e;
            10'd162:  Instruction <= 32'h24090001;
            10'd163:  Instruction <= 32'h10c9001e;
            10'd164:  Instruction <= 32'h24090002;
            10'd165:  Instruction <= 32'h10c9001e;
            10'd166:  Instruction <= 32'h24090003;
            10'd167:  Instruction <= 32'h10c9001e;
            10'd168:  Instruction <= 32'h24090004;
            10'd169:  Instruction <= 32'h10c9001e;
            10'd170:  Instruction <= 32'h24090005;
            10'd171:  Instruction <= 32'h10c9001e;
            10'd172:  Instruction <= 32'h24090006;
            10'd173:  Instruction <= 32'h10c9001e;
            10'd174:  Instruction <= 32'h24090007;
            10'd175:  Instruction <= 32'h10c9001e;
            10'd176:  Instruction <= 32'h24090008;
            10'd177:  Instruction <= 32'h10c9001e;
            10'd178:  Instruction <= 32'h24090009;
            10'd179:  Instruction <= 32'h10c9001e;
            10'd180:  Instruction <= 32'h2409000a;
            10'd181:  Instruction <= 32'h10c9001e;
            10'd182:  Instruction <= 32'h2409000b;
            10'd183:  Instruction <= 32'h10c9001e;
            10'd184:  Instruction <= 32'h2409000c;
            10'd185:  Instruction <= 32'h10c9001e;
            10'd186:  Instruction <= 32'h2409000d;
            10'd187:  Instruction <= 32'h10c9001e;
            10'd188:  Instruction <= 32'h2409000e;
            10'd189:  Instruction <= 32'h10c9001e;
            10'd190:  Instruction <= 32'h2409000f;
            10'd191:  Instruction <= 32'h10c9001e;
            10'd192:  Instruction <= 32'h24060040;
            10'd193:  Instruction <= 32'h081000e0;
            10'd194:  Instruction <= 32'h24060079;
            10'd195:  Instruction <= 32'h081000e0;
            10'd196:  Instruction <= 32'h24060024;
            10'd197:  Instruction <= 32'h081000e0;
            10'd198:  Instruction <= 32'h24060030;
            10'd199:  Instruction <= 32'h081000e0;
            10'd200:  Instruction <= 32'h24060019;
            10'd201:  Instruction <= 32'h081000e0;
            10'd202:  Instruction <= 32'h24060012;
            10'd203:  Instruction <= 32'h081000e0;
            10'd204:  Instruction <= 32'h24060002;
            10'd205:  Instruction <= 32'h081000e0;
            10'd206:  Instruction <= 32'h24060078;
            10'd207:  Instruction <= 32'h081000e0;
            10'd208:  Instruction <= 32'h24060000;
            10'd209:  Instruction <= 32'h081000e0;
            10'd210:  Instruction <= 32'h24060010;
            10'd211:  Instruction <= 32'h081000e0;
            10'd212:  Instruction <= 32'h24060008;
            10'd213:  Instruction <= 32'h081000e0;
            10'd214:  Instruction <= 32'h24060003;
            10'd215:  Instruction <= 32'h081000e0;
            10'd216:  Instruction <= 32'h24060046;
            10'd217:  Instruction <= 32'h081000e0;
            10'd218:  Instruction <= 32'h24060021;
            10'd219:  Instruction <= 32'h081000e0;
            10'd220:  Instruction <= 32'h24060006;
            10'd221:  Instruction <= 32'h081000e0;
            10'd222:  Instruction <= 32'h2406000e;
            10'd223:  Instruction <= 32'h081000e0;
            10'd224:  Instruction <= 32'h20c60b00;
            10'd225:  Instruction <= 32'h00083c00;
            10'd226:  Instruction <= 32'h00073c02;
            10'd227:  Instruction <= 32'h00073b02;
            10'd228:  Instruction <= 32'h24090000;
            10'd229:  Instruction <= 32'h10e9001e;
            10'd230:  Instruction <= 32'h24090001;
            10'd231:  Instruction <= 32'h10e9001e;
            10'd232:  Instruction <= 32'h24090002;
            10'd233:  Instruction <= 32'h10e9001e;
            10'd234:  Instruction <= 32'h24090003;
            10'd235:  Instruction <= 32'h10e9001e;
            10'd236:  Instruction <= 32'h24090004;
            10'd237:  Instruction <= 32'h10e9001e;
            10'd238:  Instruction <= 32'h24090005;
            10'd239:  Instruction <= 32'h10e9001e;
            10'd240:  Instruction <= 32'h24090006;
            10'd241:  Instruction <= 32'h10e9001e;
            10'd242:  Instruction <= 32'h24090007;
            10'd243:  Instruction <= 32'h10e9001e;
            10'd244:  Instruction <= 32'h24090008;
            10'd245:  Instruction <= 32'h10e9001e;
            10'd246:  Instruction <= 32'h24090009;
            10'd247:  Instruction <= 32'h10e9001e;
            10'd248:  Instruction <= 32'h2409000a;
            10'd249:  Instruction <= 32'h10e9001e;
            10'd250:  Instruction <= 32'h2409000b;
            10'd251:  Instruction <= 32'h10e9001e;
            10'd252:  Instruction <= 32'h2409000c;
            10'd253:  Instruction <= 32'h10e9001e;
            10'd254:  Instruction <= 32'h2409000d;
            10'd255:  Instruction <= 32'h10e9001e;
            10'd256:  Instruction <= 32'h2409000e;
            10'd257:  Instruction <= 32'h10e9001e;
            10'd258:  Instruction <= 32'h2409000f;
            10'd259:  Instruction <= 32'h10e9001e;
            10'd260:  Instruction <= 32'h24070040;
            10'd261:  Instruction <= 32'h08100124;
            10'd262:  Instruction <= 32'h24070079;
            10'd263:  Instruction <= 32'h08100124;
            10'd264:  Instruction <= 32'h24070024;
            10'd265:  Instruction <= 32'h08100124;
            10'd266:  Instruction <= 32'h24070030;
            10'd267:  Instruction <= 32'h08100124;
            10'd268:  Instruction <= 32'h24070019;
            10'd269:  Instruction <= 32'h08100124;
            10'd270:  Instruction <= 32'h24070012;
            10'd271:  Instruction <= 32'h08100124;
            10'd272:  Instruction <= 32'h24070002;
            10'd273:  Instruction <= 32'h08100124;
            10'd274:  Instruction <= 32'h24070078;
            10'd275:  Instruction <= 32'h08100124;
            10'd276:  Instruction <= 32'h24070000;
            10'd277:  Instruction <= 32'h08100124;
            10'd278:  Instruction <= 32'h24070010;
            10'd279:  Instruction <= 32'h08100124;
            10'd280:  Instruction <= 32'h24070008;
            10'd281:  Instruction <= 32'h08100124;
            10'd282:  Instruction <= 32'h24070003;
            10'd283:  Instruction <= 32'h08100124;
            10'd284:  Instruction <= 32'h24070046;
            10'd285:  Instruction <= 32'h08100124;
            10'd286:  Instruction <= 32'h24070021;
            10'd287:  Instruction <= 32'h08100124;
            10'd288:  Instruction <= 32'h24070006;
            10'd289:  Instruction <= 32'h08100124;
            10'd290:  Instruction <= 32'h2407000e;
            10'd291:  Instruction <= 32'h08100124;
            10'd292:  Instruction <= 32'h20e70700;
            10'd293:  Instruction <= 32'h24080000;
            10'd294:  Instruction <= 32'h240903e8;
            10'd295:  Instruction <= 32'h200407a4;
            10'd296:  Instruction <= 32'hae840000;
            10'd297:  Instruction <= 32'h21080001;
            10'd298:  Instruction <= 32'h0109082a;
            10'd299:  Instruction <= 32'h1420fffb;
            10'd300:  Instruction <= 32'h24080000;
            10'd301:  Instruction <= 32'h240903e8;
            10'd302:  Instruction <= 32'h20050ec0;
            10'd303:  Instruction <= 32'hae850000;
            10'd304:  Instruction <= 32'h21080001;
            10'd305:  Instruction <= 32'h0109082a;
            10'd306:  Instruction <= 32'h1420fffb;
            10'd307:  Instruction <= 32'h24080000;
            10'd308:  Instruction <= 32'h240903e8;
            10'd309:  Instruction <= 32'h20060dc0;
            10'd310:  Instruction <= 32'hae860000;
            10'd311:  Instruction <= 32'h21080001;
            10'd312:  Instruction <= 32'h0109082a;
            10'd313:  Instruction <= 32'h1420fffb;
            10'd314:  Instruction <= 32'h24080000;
            10'd315:  Instruction <= 32'h240903e8;
            10'd316:  Instruction <= 32'h20070ba4;
            10'd317:  Instruction <= 32'hae870000;
            10'd318:  Instruction <= 32'h21080001;
            10'd319:  Instruction <= 32'h0109082a;
            10'd320:  Instruction <= 32'h1420fffb;
            10'd321:  Instruction <= 32'h08100125;
            10'd322:  Instruction <= 32'h24121068;
            10'd323:  Instruction <= 32'h24080000;
            10'd324:  Instruction <= 32'hae480000;
            10'd325:  Instruction <= 32'h24080001;
            10'd326:  Instruction <= 32'h240affff;
            10'd327:  Instruction <= 32'h00124821;
            10'd328:  Instruction <= 32'h22490004;
            10'd329:  Instruction <= 32'had2a0000;
            10'd330:  Instruction <= 32'h21290004;
            10'd331:  Instruction <= 32'h21080001;
            10'd332:  Instruction <= 32'h0110082a;
            10'd333:  Instruction <= 32'h1420fffb;
            10'd334:  Instruction <= 32'h24080001;
            10'd335:  Instruction <= 32'h24090000;
            10'd336:  Instruction <= 32'h240a0000;
            10'd337:  Instruction <= 32'h00095940;
            10'd338:  Instruction <= 32'h016a5820;
            10'd339:  Instruction <= 32'h000b5880;
            10'd340:  Instruction <= 32'h00ab6020;
            10'd341:  Instruction <= 32'h8d8d0000;
            10'd342:  Instruction <= 32'h2001ffff;
            10'd343:  Instruction <= 32'h102d000f;
            10'd344:  Instruction <= 32'h00099880;
            10'd345:  Instruction <= 32'h02536020;
            10'd346:  Instruction <= 32'h8d8e0000;
            10'd347:  Instruction <= 32'h2001ffff;
            10'd348:  Instruction <= 32'h102e000a;
            10'd349:  Instruction <= 32'h000a9880;
            10'd350:  Instruction <= 32'h02536020;
            10'd351:  Instruction <= 32'h8d8f0000;
            10'd352:  Instruction <= 32'h01cda020;
            10'd353:  Instruction <= 32'h2001ffff;
            10'd354:  Instruction <= 32'h102f0003;
            10'd355:  Instruction <= 32'h028f082a;
            10'd356:  Instruction <= 32'h14200001;
            10'd357:  Instruction <= 32'h08100167;
            10'd358:  Instruction <= 32'had940000;
            10'd359:  Instruction <= 32'h214a0001;
            10'd360:  Instruction <= 32'h0150082a;
            10'd361:  Instruction <= 32'h1420ffe7;
            10'd362:  Instruction <= 32'h21290001;
            10'd363:  Instruction <= 32'h0130082a;
            10'd364:  Instruction <= 32'h1420ffe3;
            10'd365:  Instruction <= 32'h21080001;
            10'd366:  Instruction <= 32'h0110082a;
            10'd367:  Instruction <= 32'h1420ffdf;
            10'd368:  Instruction <= 32'h24080008;
            10'd369:  Instruction <= 32'hae480004;
            10'd370:  Instruction <= 32'h24080003;
            10'd371:  Instruction <= 32'hae480008;
            10'd372:  Instruction <= 32'h24080005;
            10'd373:  Instruction <= 32'hae48000c;
            10'd374:  Instruction <= 32'h2408000a;
            10'd375:  Instruction <= 32'hae480010;
            10'd376:  Instruction <= 32'h24080008;
            10'd377:  Instruction <= 32'hae480014;
            10'd378:  Instruction <= 32'h03e00008;




			// -------- Paste Binary Instruction Above
			
			default: Instruction <= 32'h00000000;
		endcase
		
endmodule
